module mem_ram #(
    parameter WIDTH = 8
) (
    
);
    
endmodule